library IEEE;
use IEEE.std_logic_1164.all;

entity ent is
port (d : in std_logic_vector(3 downto 0);
			clk, load, shift : in std_logic;
			qout : out std_logic);
end ent;

architecture arch of ent is

    

begin

end arch ; -- arch